module bin2bcd #(
  parameter WIDTH = 8
)(
  input logic   x,
  output logic  bcd
);

always_ff @ (posedge clk)



endmodule
